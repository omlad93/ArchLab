module main;
  // FILL HERE
endmodule

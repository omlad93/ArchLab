module halfadder(a,b,sum,carry);
  input a,b;
  output sum, carry;
  wire sum, carry;

  xor g0(/* FILL HERE */);
  and g1(/* FILL HERE */);
endmodule

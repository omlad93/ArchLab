module parity(clk, in, reset, out);

   input clk, in, reset;
   output out;

   reg 	  out;
   reg 	  state;

   localparam zero=0, one=1;

   always @(posedge clk)
     begin
	if (reset)
	  state <= zero;
	else
	  case (state)
	    // FILL HERE
	  endcase
     end

   always @(state) 
     begin
	case (state)
	    // FILL HERE
	endcase
     end

endmodule

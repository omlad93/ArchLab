module fulladder( sum, co, a, b, ci);

  input   a, b, ci;
  output  sum, co;

  // FILL HERE

endmodule
